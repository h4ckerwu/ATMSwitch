package virtual_interfaces;

    typedef virtual Utopia vUtopia;
    typedef virtual Utopia.TB_Rx vUtopiaRx;
    typedef virtual Utopia.TB_Tx vUtopiaTx;

    typedef virtual cpu_ifc vCPU;
    typedef virtual cpu_ifc.Test vCPU_T;

endpackage

